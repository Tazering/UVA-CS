-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
-- CREATED		"Sat Sep 10 21:22:33 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY majority_voter0 IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		Z :  OUT  STD_LOGIC
	);
END majority_voter0;

ARCHITECTURE bdf_type OF majority_voter0 IS 

SIGNAL	wire0 :  STD_LOGIC;
SIGNAL	wire1 :  STD_LOGIC;
SIGNAL	wire2 :  STD_LOGIC;


BEGIN 



wire0 <= A AND B;


wire1 <= B AND C;


wire2 <= C AND A;


Z <= wire1 OR wire2 OR wire0;


END bdf_type;